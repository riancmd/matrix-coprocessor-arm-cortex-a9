module opp_M()

endmodule