module alu3(input [600:00] a); 
	
endmodule